`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
module G_function(clk, W4, g_out, rc_in);
 input clk;
 input [31:0] W4;
 input [7:0] rc_in;
 output [31:0] g_out;
 reg [7:0] LUT[0:15][0:15];
 reg [7:0] v0, v1, v2, v3; 
   
 initial begin
 LUT[0][0] <= 8'h63; 
 LUT[0][1] <= 8'h7C; 
 LUT[0][2] <= 8'h77;
 LUT[0][3] <= 8'h7B; 
 LUT[0][4] <= 8'hF2;
 LUT[0][5] <= 8'h6B; 
 LUT[0][6] <= 8'h6F; 
 LUT[0][7] <= 8'hC5;
 LUT[0][8] <= 8'h30; 
 LUT[0][9] <= 8'h01;
 LUT[0][10] <= 8'h67;
 LUT[0][11] <= 8'h2B;
 LUT[0][12] <= 8'hFE;
 LUT[0][13] <= 8'hD7;
 LUT[0][14] <= 8'hAB; 
 LUT[0][15] <= 8'h76;
 LUT[1][0] <= 8'hCA;
 LUT[1][1] <= 8'h82; 
 LUT[1][2] <= 8'hC9;
 LUT[1][3] <= 8'h7D; 
 LUT[1][4] <= 8'hFA;
 LUT[1][5] <= 8'h59;
 LUT[1][6] <= 8'h47;
 LUT[1][7] <= 8'hF0;
 LUT[1][8] <= 8'hAD;
 LUT[1][9] <= 8'hD4;
 LUT[1][10] <= 8'hA2;
 LUT[1][11] <= 8'hAF;
 LUT[1][12] <= 8'h9C;
 LUT[1][13] <= 8'hA4;
 LUT[1][14] <= 8'h72;
 LUT[1][15] <= 8'hC0;
 LUT[2][0] <= 8'hB7;
 LUT[2][1] <= 8'hFD;
 LUT[2][2] <= 8'h93;
 LUT[2][3] <= 8'h26;
 LUT[2][4] <= 8'h36;
 LUT[2][5] <= 8'h3F;
 LUT[2][6] <= 8'hF7;
 LUT[2][7] <= 8'hCC;
 LUT[2][8] <= 8'h34;
 LUT[2][9] <= 8'hA5;
 LUT[2][10] <= 8'hE5;
 LUT[2][11] <= 8'hF1;
 LUT[2][12] <= 8'h71;
 LUT[2][13] <= 8'hD8; 
 LUT[2][14] <= 8'h31;
 LUT[2][15] <= 8'h15;
 LUT[3][0] <= 8'h04; 
 LUT[3][1] <= 8'hC7; 
 LUT[3][2] <= 8'h23;
 LUT[3][3] <= 8'hC3;
 LUT[3][4] <= 8'h18; 
 LUT[3][5] <= 8'h96;
 LUT[3][6] <= 8'h05; 
 LUT[3][7] <= 8'h9A;
 LUT[3][8] <= 8'h07; 
 LUT[3][9] <= 8'h12;
 LUT[3][10] <= 8'h80;
 LUT[3][11] <= 8'hE2;
 LUT[3][12] <= 8'hEB;
 LUT[3][13] <= 8'h27;
 LUT[3][14] <= 8'hB2;
 LUT[3][15] <= 8'h75;
 LUT[4][0] <= 8'h09; 
 LUT[4][1] <= 8'h83;
 LUT[4][2] <= 8'h2C; 
 LUT[4][3] <= 8'h1A; 
 LUT[4][4] <= 8'h1B;
 LUT[4][5] <= 8'h6E; 
 LUT[4][6] <= 8'h5A; 
 LUT[4][7] <= 8'hA0;
 LUT[4][8] <= 8'h52; 
 LUT[4][9] <= 8'h3B; 
 LUT[4][10] <= 8'hD6;
 LUT[4][11] <= 8'hB3; 
 LUT[4][12] <= 8'h29;
 LUT[4][13] <= 8'hE3;
 LUT[4][14] <= 8'h2F;
 LUT[4][15] <= 8'h84;
 LUT[5][0] <= 8'h53;
 LUT[5][1] <= 8'hD1; 
 LUT[5][2] <= 8'h00; 
 LUT[5][3] <= 8'hED;
 LUT[5][4] <= 8'h20; 
 LUT[5][5] <= 8'hFC;
 LUT[5][6] <= 8'hB1; 
 LUT[5][7] <= 8'h5B;
 LUT[5][8] <= 8'h6A; 
 LUT[5][9] <= 8'hCB; 
 LUT[5][10] <= 8'hBE; 
 LUT[5][11] <= 8'h39; 
 LUT[5][12] <= 8'h4A;
 LUT[5][13] <= 8'h4C;
 LUT[5][14] <= 8'h58; 
 LUT[5][15] <= 8'hCF;
 LUT[6][0] <= 8'hD0;
LUT[6][1] <= 8'hEF; 
LUT[6][2] <= 8'hAA;
LUT[6][3] <= 8'hFB; 
LUT[6][4] <= 8'h43; 
LUT[6][5] <= 8'h4D; 
LUT[6][6] <= 8'h33;
LUT[6][7] <= 8'h85; 
LUT[6][8] <= 8'h45; 
LUT[6][9] <= 8'hF9;
LUT[6][10] <= 8'h02;
LUT[6][11] <= 8'h7F;
LUT[6][12] <= 8'h50;
LUT[6][13] <= 8'h3C;
LUT[6][14] <= 8'h9F;
LUT[6][15] <= 8'hA8;
LUT[7][0] <= 8'h51;
LUT[7][1] <= 8'hA3;
LUT[7][2] <= 8'h40; 
LUT[7][3] <= 8'h8F; 
LUT[7][4] <= 8'h92;
LUT[7][5] <= 8'h9D;  
LUT[7][6] <= 8'h38;
LUT[7][7] <= 8'hF5;
LUT[7][8] <= 8'hBC;
LUT[7][9] <= 8'hB6;
LUT[7][10] <= 8'hDA;
LUT[7][11] <= 8'h21; 
LUT[7][12] <= 8'h10;
LUT[7][13] <= 8'hFF;
LUT[7][14] <= 8'hF3;
LUT[7][15] <= 8'hD2;
LUT[8][0] <= 8'hCD;
LUT[8][1] <= 8'h0C; 
LUT[8][2] <= 8'h13; 
LUT[8][3] <= 8'hEC;
LUT[8][4] <= 8'h5F;
LUT[8][5] <= 8'h97;
LUT[8][6] <= 8'h44; 
LUT[8][7] <= 8'h17; 
LUT[8][8] <= 8'hC4;
LUT[8][9] <= 8'hA7; 
LUT[8][10] <= 8'h7E; 
LUT[8][11] <= 8'h3D; 
LUT[8][12] <= 8'h64; 
LUT[8][13] <= 8'h5D; 
LUT[8][14] <= 8'h19;  
LUT[8][15] <= 8'h73;
LUT[9][0] <= 8'h60; 
LUT[9][1] <= 8'h81; 
LUT[9][2] <= 8'h4F; 
LUT[9][3] <= 8'hDC;
LUT[9][4] <= 8'h22;  
LUT[9][5] <= 8'h2A;
LUT[9][6] <= 8'h90; 
LUT[9][7] <= 8'h88; 
LUT[9][8] <= 8'h46; 
LUT[9][9] <= 8'hEE;
LUT[9][10] <= 8'hB8;
LUT[9][11] <= 8'h14; 
LUT[9][12] <= 8'hDE;
LUT[9][13] <= 8'h5E; 
LUT[9][14] <= 8'h0B; 
LUT[9][15] <= 8'hDB;
LUT[10][0] <= 8'hE0;
LUT[10][1] <= 8'h32; 
LUT[10][2] <= 8'h3A;
LUT[10][3] <= 8'h0A; 
LUT[10][4] <= 8'h49;
LUT[10][5] <= 8'h06;  
LUT[10][6] <= 8'h24; 
LUT[10][7] <= 8'h5C; 
LUT[10][8] <= 8'hC2;
LUT[10][9] <= 8'hD3;  
LUT[10][10] <= 8'hAC;  
LUT[10][11] <= 8'h62;
LUT[10][12] <= 8'h91; 
LUT[10][13] <= 8'h95;  
LUT[10][14] <= 8'hE4; 
LUT[10][15] <= 8'h79; 
LUT[11][0] <= 8'hE7; 
LUT[11][1] <= 8'hC8; 
LUT[11][2] <= 8'h37;  
LUT[11][3] <= 8'h6D;
LUT[11][4] <= 8'h8D;  
LUT[11][5] <= 8'hD5;  
LUT[11][6] <= 8'h4E;  
LUT[11][7] <= 8'hA9;  
LUT[11][8] <= 8'h6C; 
LUT[11][9] <= 8'h56;  
LUT[11][10] <= 8'hF4;    
LUT[11][11] <= 8'hEA;  
LUT[11][12] <= 8'h65; 
LUT[11][13] <= 8'h7A; 
LUT[11][14] <= 8'hAE; 
LUT[11][15] <= 8'h08;
LUT[12][0] <= 8'hBA;  
LUT[12][1] <= 8'h78; 
LUT[12][2] <= 8'h25;  
LUT[12][3] <= 8'h2E; 
LUT[12][4] <= 8'h1C;  
LUT[12][5] <= 8'hA6;  
LUT[12][6] <= 8'hB4; 
LUT[12][7] <= 8'hC6; 
LUT[12][8] <= 8'hE8;
LUT[12][9] <= 8'hDD; 
LUT[12][10] <= 8'h74; 
LUT[12][11] <= 8'h1F;   
LUT[12][12] <= 8'h4B; 
LUT[12][13] <= 8'hBD;  
LUT[12][14] <= 8'h8B; 
LUT[12][15] <= 8'h8A;
LUT[13][0] <= 8'h70;
LUT[13][1] <= 8'h3E; 
LUT[13][2] <= 8'hB5; 
LUT[13][3] <= 8'h66;  
LUT[13][4] <= 8'h48; 
LUT[13][5] <= 8'h03; 
LUT[13][6] <= 8'hF6;
LUT[13][7] <= 8'h0E;  
LUT[13][8] <= 8'h61;  
LUT[13][9] <= 8'h35; 
LUT[13][10] <= 8'h57;
LUT[13][11] <= 8'hB9; 
LUT[13][12] <= 8'h86;
LUT[13][13] <= 8'hC1;  
LUT[13][14] <= 8'h1D; 
LUT[13][15] <= 8'h9E;
LUT[14][0] <= 8'hE1; 
LUT[14][1] <= 8'hF8;
LUT[14][2] <= 8'h98; 
LUT[14][3] <= 8'h11; 
LUT[14][4] <= 8'h69;  
LUT[14][5] <= 8'hD9; 
LUT[14][6] <= 8'h8E; 
LUT[14][7] <= 8'h94;
LUT[14][8] <= 8'h9B; 
LUT[14][9] <= 8'h1E; 
LUT[14][10] <= 8'h87; 
LUT[14][11] <= 8'hE9; 
LUT[14][12] <= 8'hCE;   
LUT[14][13] <= 8'h55;  
LUT[14][14] <= 8'h28;  
LUT[14][15] <= 8'hDF;
LUT[15][0] <= 8'h8C; 
LUT[15][1] <= 8'hA1;  
LUT[15][2] <= 8'h89; 
LUT[15][3] <= 8'h0D;  
LUT[15][4] <= 8'hBF;  
LUT[15][5] <= 8'hE6;  
LUT[15][6] <= 8'h42;  
LUT[15][7] <= 8'h68;  
LUT[15][8] <= 8'h41;   
LUT[15][9] <= 8'h99;  
LUT[15][10] <= 8'h2D; 
LUT[15][11] <= 8'h0F;  
LUT[15][12] <= 8'hB0; 
LUT[15][13] <= 8'h54;  
LUT[15][14] <= 8'hBB;  
LUT[15][15] <= 8'h16;
end

always@(posedge clk)
begin
v0 <= W4[31:24];
v1 <= W4[23:16];
v2 <= W4[15:8];
v3 <= W4[7:0];
end

assign g_out[31:24] = rc_in + LUT[v1[7:4]][v1[3:0]];
assign g_out[23:16] = LUT[v2[7:4]][v2[3:0]];
assign g_out[15:8] = LUT[v3[7:4]][v3[3:0]];
assign g_out[7:0] = LUT[v0[7:4]][v0[3:0]]; 

endmodule
